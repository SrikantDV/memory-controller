interface power_intf();

endinterface

module mc_timing();
and
or
nand
nor();
endmodule

DFT, Physical Design will be done on this wrong netlist
STA
Layout done on wrong netlist
Chip will be manufactured with a wrong netlist

//rtl file list
`include "mc_adr_sel.v"
`include "mc_cs_rf.v"
`include "mc_defines.v"
`include "mc_dp.v"
`include "mc_incn_r.v"
`include "mc_mem_if.v"
`include "mc_obct.v"
`include "mc_obct_top.v"
`include "mc_rd_fifo.v"
`include "mc_refresh.v"
`include "mc_rf.v"
`include "mc_timing.v"
`include "mc_top.v"
`include "mc_wb_if.v"
`include "timescale.v"

//testbench files
`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "mc_common.sv"
`include "wb_tx.sv"
`include "mem_intf.sv"
`include "wb_interface.sv"

`include "wb_seq_lib.sv"
`include "wb_monitor.sv"
`include "wb_coverage.sv"
`include "wb_sqr.sv"
`include "wb_driver.sv"
`include "wb_agent.sv"
`include "mc_env.sv"
`include "mc_test_lib.sv"
`include "mem_top.sv"
